`timescale 1ns / 1ps

module draw_track
#(parameter
    RECT_WIDTH = 16,
    RECT_LENGTH = 16,
    ADDR_WIDTH = 16
)
(
    input wire [10:0] hcount_in,
    input wire hsync_in,
    input wire hblnk_in,
    input wire [10:0] vcount_in,
    input wire vsync_in,
    input wire vblnk_in,
    input wire pclk,
    input wire rst,
    input wire visible,
    input wire [11:0] rgb_in,
    input wire [11:0] rgb_pixel,
    output reg [10:0] hcount_out,
    output reg hsync_out,
    output reg hblnk_out,
    output reg [10:0] vcount_out,
    output reg vsync_out,
    output reg vblnk_out,
    output reg [11:0] rgb_out,
    output reg [ADDR_WIDTH-1:0] pixel_addr
);

localparam SCREEN_WIDTH = 1024;
localparam SCREEN_HEIGHT = 768;

reg [11:0] rgb_out_nxt;
wire [10:0] xpos, ypos, xpos_nxt, ypos_nxt;
reg [10:0] tile_x_pos, tile_y_pos;
reg [ADDR_WIDTH-1:0] pixel_addr_nxt;
reg [10:0] addrx, addry;
wire [10:0] vcount_delayed, hcount_delayed;
wire hsync_delayed, vsync_delayed, hblnk_delayed, vblnk_delayed;

assign xpos = (hcount_in / 16);
assign ypos = (vcount_in / 16);

always @(posedge pclk)
    if(rst)
    begin
        hcount_out <= 0;
        hsync_out <= 0;
        hblnk_out <= 0;
        vcount_out <= 0;
        vsync_out <= 0;
        vblnk_out <= 0;
        rgb_out <= 0;
        pixel_addr <= 0;
    end
    else
    begin
        hcount_out <= hcount_delayed;
        hsync_out <= hsync_delayed;
        hblnk_out <= hblnk_delayed;
        vcount_out <= vcount_delayed;
        vsync_out <= vsync_delayed;
        vblnk_out <= vblnk_delayed;
        rgb_out <= rgb_out_nxt;
        pixel_addr <= pixel_addr_nxt;
    end

always @*
begin
    addrx = hcount_in + tile_x_pos - (xpos * 16);
    addry = vcount_in + tile_y_pos - (ypos * 16);
    rgb_out_nxt = rgb_in;
    pixel_addr_nxt = 0;
    if(visible)
    begin
        if(hcount_in >= 0 && hcount_in < (SCREEN_WIDTH) && vcount_in >= 0 && vcount_in < (SCREEN_HEIGHT))
        begin
            rgb_out_nxt = rgb_pixel;
            pixel_addr_nxt = { (addry[(ADDR_WIDTH/2)-1:0]), (addrx[(ADDR_WIDTH/2)-1:0]) };
        end
    end
end

always @*
case ((ypos * 64) + xpos)
    0:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    4:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    5:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    6:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    7:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    8:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    9:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    10:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    11:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    12:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    13:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    14:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    15:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    16:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    17:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    18:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    19:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    20:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    21:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    22:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    23:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    24:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    25:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    26:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    27:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    28:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    29:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    30:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    31:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    32:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    33:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    34:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    35:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    36:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    37:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    38:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    39:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    40:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    41:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    42:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    43:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    44:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    45:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    46:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    47:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    48:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    49:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    50:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    51:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    52:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    53:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    54:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    55:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    56:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    57:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    58:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    59:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    60:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    61:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    62:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    63:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    64:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    65:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    66:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    67:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    68:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    69:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    70:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    71:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    72:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    73:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    74:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    75:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    76:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    77:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    78:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    79:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    80:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    81:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    82:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    83:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    84:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    85:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    86:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    87:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    88:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    89:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    90:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    91:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    92:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    93:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    94:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    95:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    96:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    97:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    98:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    99:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    100:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    101:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    102:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    103:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    104:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    105:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    106:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    107:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    108:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    109:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    110:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    111:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    112:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    113:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    114:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    115:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    116:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    117:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    118:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    119:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    120:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    121:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    122:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    123:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    124:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    125:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    126:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    127:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    128:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    129:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    130:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    131:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    132:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    133:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    134:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    135:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    136:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    137:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    138:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    139:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    140:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    141:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    142:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    143:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    144:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    145:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    146:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    147:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    148:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    149:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    150:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    151:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    152:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    153:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    154:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    155:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    156:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    157:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    158:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    159:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    160:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    161:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    162:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    163:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    164:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    165:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    166:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    167:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    168:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    169:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    170:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    171:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    172:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    173:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    174:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    175:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    176:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    177:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    178:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    179:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    180:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    181:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    182:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    183:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    184:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    185:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    186:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    187:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    188:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    189:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    190:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    191:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    192:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    193:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    194:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    195:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    196:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    197:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    198:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    199:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    200:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    201:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    202:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    203:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    204:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    205:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    206:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    207:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    208:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    209:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    210:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    211:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    212:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    213:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    214:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    215:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    216:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    217:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    218:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    219:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    220:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    221:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    222:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    223:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    224:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    225:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    226:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    227:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    228:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    229:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    230:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    231:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    232:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    233:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    234:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    235:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    236:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    237:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    238:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    239:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    240:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    241:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    242:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    243:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    244:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    245:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    246:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    247:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    248:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    249:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    250:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    251:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    252:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    253:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    254:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    255:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    256:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    257:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    258:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    259:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    260:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    261:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    262:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    263:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    264:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    265:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    266:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    267:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    268:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    269:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    270:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    271:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    272:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    273:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    274:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    275:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    276:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    277:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    278:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    279:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    280:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    281:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    282:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    283:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    284:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    285:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    286:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    287:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    288:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    289:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    290:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    291:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    292:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    293:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    294:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    295:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    296:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    297:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    298:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    299:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    300:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    301:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    302:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    303:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    304:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    305:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    306:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    307:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    308:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    309:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    310:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    311:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    312:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    313:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    314:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    315:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    316:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    317:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    318:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    319:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    320:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    321:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    322:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    323:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    324:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    325:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    326:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    327:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    328:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    329:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    330:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    331:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    332:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    333:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    334:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    335:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    336:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    337:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    338:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    339:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    340:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    341:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    342:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    343:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    344:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    345:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    346:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    347:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    348:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    349:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    350:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    351:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    352:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    353:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    354:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    355:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    356:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    357:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    358:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    359:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    360:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    361:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    362:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    363:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    364:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    365:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    366:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    367:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    368:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    369:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    370:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    371:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    372:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    373:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    374:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    375:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    376:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    377:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    378:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    379:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    380:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    381:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    382:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    383:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    384:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    385:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    386:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    387:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    388:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    389:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    390:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    391:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    392:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    393:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    394:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    395:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    396:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    397:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    398:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    399:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    400:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    401:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    402:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    403:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    404:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    405:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    406:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    407:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    408:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    409:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    410:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    411:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    412:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    413:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    414:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    415:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    416:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    417:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    418:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    419:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    420:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    421:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    422:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    423:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    424:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    425:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    426:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    427:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    428:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    429:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    430:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    431:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    432:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    433:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    434:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    435:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    436:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    437:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    438:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    439:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    440:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    441:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    442:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    443:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    444:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    445:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    446:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    447:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    448:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    449:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    450:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    451:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    452:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    453:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    454:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    455:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    456:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    457:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    458:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    459:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    460:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    461:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    462:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    463:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    464:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    465:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    466:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    467:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    468:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    469:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    470:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    471:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    472:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    473:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    474:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    475:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    476:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    477:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    478:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    479:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    480:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    481:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    482:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    483:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    484:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    485:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    486:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    487:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    488:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    489:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    490:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    491:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    492:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    493:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    494:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    495:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    496:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    497:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    498:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    499:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    500:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    501:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    502:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    503:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    504:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    505:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    506:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    507:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    508:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    509:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    510:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    511:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    512:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    513:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    514:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    515:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    516:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    517:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    518:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    519:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    520:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    521:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    522:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    523:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    524:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    525:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    526:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    527:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    528:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    529:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    530:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    531:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    532:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    533:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    534:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    535:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    536:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    537:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    538:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    539:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    540:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    541:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    542:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    543:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    544:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    545:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    546:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    547:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    548:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    549:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    550:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    551:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    552:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    553:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    554:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    555:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    556:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    557:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    558:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    559:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    560:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    561:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    562:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    563:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    564:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    565:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    566:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    567:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    568:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    569:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    570:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    571:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    572:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    573:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    574:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    575:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    576:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    577:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    578:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    579:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    580:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    581:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    582:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    583:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    584:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    585:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    586:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    587:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    588:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    589:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    590:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    591:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    592:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    593:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    594:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    595:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    596:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    597:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    598:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    599:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    600:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    601:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    602:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    603:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    604:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    605:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    606:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    607:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    608:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    609:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    610:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    611:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    612:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    613:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    614:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    615:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    616:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    617:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    618:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    619:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    620:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    621:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    622:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    623:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    624:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    625:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    626:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    627:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    628:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    629:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    630:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    631:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    632:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    633:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    634:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    635:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    636:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    637:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    638:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    639:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    640:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    641:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    642:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    643:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    644:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    645:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    646:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    647:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    648:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    649:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    650:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    651:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    652:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    653:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    654:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    655:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    656:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    657:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    658:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    659:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    660:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    661:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    662:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    663:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    664:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    665:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    666:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    667:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    668:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    669:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    670:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    671:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    672:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    673:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    674:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    675:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    676:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    677:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    678:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    679:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    680:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    681:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    682:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    683:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    684:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    685:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    686:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    687:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    688:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    689:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    690:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    691:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    692:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    693:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    694:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    695:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    696:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    697:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    698:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    699:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    700:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    701:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    702:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    703:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    704:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    705:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    706:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    707:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    708:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    709:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    710:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    711:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    712:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    713:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    714:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    715:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    716:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    717:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    718:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    719:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    720:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    721:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    722:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    723:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    724:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    725:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    726:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    727:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    728:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    729:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    730:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    731:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    732:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    733:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    734:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    735:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    736:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    737:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    738:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    739:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    740:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    741:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    742:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    743:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    744:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    745:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    746:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    747:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    748:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    749:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    750:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    751:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    752:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    753:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    754:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    755:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    756:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    757:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    758:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    759:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    760:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    761:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    762:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    763:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    764:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    765:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    766:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    767:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    768:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    769:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    770:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    771:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    772:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    773:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    774:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    775:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    776:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    777:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    778:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    779:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    780:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    781:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    782:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    783:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    784:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    785:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    786:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    787:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    788:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    789:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    790:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    791:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    792:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    793:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    794:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    795:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    796:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    797:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    798:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    799:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    800:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    801:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    802:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    803:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    804:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    805:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    806:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    807:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    808:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    809:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    810:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    811:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    812:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    813:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    814:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    815:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    816:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    817:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    818:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    819:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    820:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    821:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    822:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    823:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    824:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    825:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    826:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    827:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    828:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    829:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    830:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    831:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    832:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    833:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    834:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    835:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    836:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    837:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    838:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    839:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    840:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    841:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    842:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    843:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    844:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    845:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    846:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    847:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    848:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    849:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    850:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    851:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    852:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    853:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    854:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    855:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    856:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    857:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    858:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    859:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    860:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    861:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    862:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    863:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    864:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    865:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    866:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    867:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    868:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    869:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    870:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    871:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    872:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    873:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    874:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    875:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    876:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    877:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    878:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    879:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    880:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    881:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    882:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    883:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    884:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    885:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    886:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    887:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    888:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    889:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    890:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    891:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    892:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    893:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    894:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    895:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    896:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    897:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    898:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    899:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    900:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    901:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    902:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    903:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    904:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    905:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    906:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    907:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    908:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    909:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    910:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    911:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    912:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    913:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    914:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    915:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    916:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    917:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    918:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    919:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    920:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    921:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    922:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    923:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    924:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    925:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    926:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    927:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    928:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    929:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    930:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    931:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    932:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    933:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    934:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    935:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    936:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    937:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    938:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    939:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    940:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    941:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    942:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    943:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    944:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    945:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    946:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    947:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    948:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    949:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    950:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    951:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    952:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    953:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    954:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    955:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    956:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    957:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    958:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    959:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    960:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    961:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    962:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    963:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    964:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    965:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    966:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    967:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    968:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    969:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    970:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    971:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    972:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    973:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    974:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    975:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    976:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    977:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    978:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    979:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    980:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    981:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    982:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    983:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    984:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    985:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    986:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    987:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    988:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    989:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    990:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    991:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    992:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    993:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    994:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    995:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    996:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    997:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    998:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    999:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1000:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1001:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1002:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1003:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1004:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1005:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1006:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1007:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1008:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1009:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1010:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1011:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1012:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1013:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1014:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1015:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1016:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1017:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1018:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1019:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1020:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1021:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1022:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1023:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1024:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1025:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1026:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1027:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1028:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1029:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1030:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1031:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1032:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1033:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1034:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1035:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1036:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1037:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1038:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1039:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1040:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1041:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1042:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1043:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1044:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1045:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1046:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1047:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1048:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1049:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1050:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1051:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1052:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1053:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1054:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1055:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1056:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1057:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1058:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1059:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1060:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1061:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1062:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1063:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1064:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1065:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1066:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1067:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1068:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1069:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1070:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1071:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1072:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1073:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1074:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1075:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1076:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1077:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1078:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1079:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1080:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1081:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1082:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1083:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1084:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1085:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1086:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1087:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1088:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1089:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1090:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1091:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1092:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1093:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1094:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1095:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1096:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1097:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1098:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1099:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1100:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1101:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1102:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1103:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1104:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1105:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1106:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1107:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1108:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1109:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1110:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1111:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1112:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1113:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1114:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1115:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1116:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1117:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1118:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1119:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1120:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1121:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1122:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1123:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1124:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1125:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1126:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1127:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1128:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1129:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1130:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1131:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1132:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1133:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1134:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1135:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1136:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1137:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1138:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1139:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1140:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1141:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1142:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1143:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1144:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1145:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1146:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1147:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1148:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1149:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1150:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1151:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1152:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1153:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1154:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1155:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1156:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1157:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1158:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1159:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1160:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1161:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1162:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1163:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1164:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1165:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1166:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1167:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1168:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1169:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1170:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1171:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1172:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1173:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1174:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1175:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1176:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1177:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1178:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1179:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1180:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1181:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1182:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1183:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1184:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1185:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1186:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1187:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1188:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1189:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1190:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1191:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1192:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1193:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1194:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1195:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1196:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1197:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1198:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1199:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1200:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1201:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1202:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1203:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1204:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1205:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1206:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1207:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1208:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1209:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1210:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1211:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1212:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1213:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1214:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1215:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1216:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1217:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1218:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1219:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1220:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1221:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1222:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1223:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1224:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1225:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1226:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1227:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1228:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1229:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1230:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1231:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1232:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1233:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1234:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1235:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1236:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1237:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1238:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1239:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1240:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1241:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1242:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1243:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1244:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1245:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1246:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1247:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1248:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1249:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1250:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1251:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1252:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1253:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1254:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1255:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1256:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1257:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1258:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1259:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1260:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1261:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1262:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1263:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1264:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1265:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1266:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1267:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1268:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1269:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1270:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1271:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1272:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1273:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1274:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1275:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1276:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1277:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1278:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1279:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1280:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1281:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1282:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1283:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1284:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1285:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1286:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1287:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1288:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1289:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1290:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1291:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1292:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1293:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1294:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1295:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1296:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1297:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1298:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1299:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1300:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1301:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1302:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1303:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1304:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1305:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1306:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1307:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1308:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1309:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1310:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1311:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1312:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1313:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1314:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1315:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1316:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1317:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1318:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1319:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1320:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1321:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1322:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1323:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1324:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1325:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1326:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1327:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1328:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1329:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1330:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1331:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1332:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1333:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1334:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1335:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1336:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1337:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1338:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1339:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1340:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1341:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1342:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1343:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1344:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1345:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1346:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1347:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1348:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1349:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1350:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1351:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1352:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1353:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1354:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1355:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1356:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1357:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1358:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1359:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1360:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1361:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1362:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1363:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1364:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1365:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1366:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1367:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1368:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1369:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1370:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1371:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1372:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1373:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1374:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1375:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1376:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1377:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1378:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1379:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1380:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1381:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1382:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1383:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1384:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1385:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1386:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1387:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1388:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1389:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1390:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1391:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1392:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1393:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1394:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1395:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1396:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1397:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1398:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1399:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1400:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1401:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1402:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1403:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1404:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1405:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1406:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1407:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1408:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1409:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1410:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1411:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1412:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1413:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1414:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1415:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1416:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1417:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1418:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1419:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1420:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1421:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1422:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1423:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1424:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1425:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1426:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1427:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1428:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1429:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1430:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1431:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1432:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1433:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1434:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1435:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1436:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1437:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1438:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1439:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1440:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1441:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1442:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1443:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1444:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1445:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1446:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1447:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1448:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1449:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1450:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1451:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1452:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1453:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1454:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1455:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1456:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1457:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1458:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1459:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1460:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1461:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1462:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1463:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1464:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1465:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1466:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1467:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1468:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1469:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1470:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1471:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1472:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1473:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1474:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1475:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1476:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1477:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1478:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1479:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1480:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1481:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1482:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1483:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1484:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1485:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1486:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1487:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1488:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1489:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1490:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1491:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1492:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1493:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1494:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1495:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1496:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1497:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1498:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1499:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1500:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1501:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1502:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1503:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1504:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1505:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1506:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1507:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1508:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1509:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1510:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1511:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1512:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1513:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1514:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1515:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1516:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1517:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1518:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1519:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1520:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1521:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1522:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1523:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1524:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1525:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1526:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1527:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1528:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1529:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1530:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1531:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1532:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1533:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1534:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1535:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1536:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1537:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1538:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1539:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1540:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1541:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1542:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1543:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1544:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1545:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1546:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1547:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1548:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1549:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1550:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1551:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1552:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1553:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1554:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1555:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1556:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1557:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1558:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1559:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1560:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1561:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1562:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1563:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1564:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1565:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1566:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1567:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1568:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1569:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1570:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1571:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1572:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1573:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1574:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1575:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1576:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1577:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1578:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1579:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1580:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1581:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1582:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1583:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1584:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1585:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1586:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1587:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1588:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1589:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1590:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1591:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1592:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1593:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1594:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1595:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1596:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1597:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1598:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1599:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1600:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1601:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1602:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1603:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1604:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1605:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1606:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1607:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1608:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1609:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1610:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1611:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1612:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1613:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1614:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1615:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1616:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1617:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1618:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1619:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1620:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1621:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1622:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1623:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1624:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1625:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1626:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1627:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1628:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1629:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1630:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1631:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1632:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1633:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1634:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1635:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1636:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1637:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1638:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1639:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1640:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1641:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1642:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1643:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1644:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1645:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1646:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1647:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1648:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1649:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1650:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1651:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1652:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1653:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1654:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1655:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1656:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1657:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1658:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1659:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1660:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1661:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1662:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1663:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1664:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1665:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1666:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1667:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1668:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1669:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1670:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1671:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1672:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1673:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1674:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1675:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1676:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1677:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1678:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1679:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1680:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1681:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1682:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1683:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1684:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1685:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1686:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1687:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1688:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1689:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1690:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1691:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1692:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1693:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1694:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1695:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1696:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1697:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1698:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1699:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1700:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1701:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1702:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1703:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 2);
    end
    1704:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1705:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1706:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1707:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1708:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1709:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1710:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1711:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1712:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1713:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1714:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1715:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1716:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1717:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1718:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1719:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1720:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1721:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1722:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1723:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1724:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1725:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1726:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1727:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1728:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1729:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1730:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1731:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1732:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1733:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1734:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1735:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1736:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1737:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1738:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1739:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1740:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1741:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1742:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1743:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1744:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1745:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1746:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 3);
    end
    1747:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1748:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1749:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1750:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1751:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1752:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1753:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1754:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1755:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1756:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1757:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1758:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1759:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1760:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1761:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1762:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1763:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1764:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1765:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1766:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1767:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1768:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1769:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1770:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1771:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1772:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1773:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1774:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1775:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1776:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1777:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1778:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1779:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1780:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1781:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1782:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1783:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1784:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1785:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1786:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1787:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1788:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1789:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1790:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1791:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1792:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1793:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1794:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1795:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1796:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1797:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1798:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1799:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1800:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1801:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1802:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1803:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1804:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1805:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1806:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1807:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1808:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1809:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1810:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1811:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1812:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1813:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1814:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1815:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1816:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1817:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1818:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1819:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1820:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1821:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1822:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1823:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1824:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1825:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1826:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1827:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1828:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1829:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1830:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1831:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1832:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1833:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1834:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1835:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1836:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1837:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1838:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1839:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1840:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1841:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1842:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1843:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1844:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1845:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1846:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1847:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1848:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1849:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1850:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1851:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1852:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1853:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1854:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1855:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1856:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1857:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1858:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1859:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1860:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1861:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1862:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1863:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1864:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1865:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1866:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1867:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1868:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1869:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1870:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1871:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1872:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1873:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1874:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1875:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1876:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1877:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1878:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1879:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1880:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1881:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1882:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1883:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1884:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1885:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1886:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1887:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1888:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1889:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1890:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1891:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1892:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1893:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1894:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1895:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1896:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1897:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1898:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1899:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1900:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1901:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1902:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1903:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1904:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1905:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1906:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1907:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1908:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1909:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1910:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1911:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1912:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1913:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1914:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1915:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1916:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1917:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1918:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1919:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1920:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1921:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1922:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1923:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1924:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1925:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1926:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1927:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1928:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 4);
    end
    1929:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1930:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1931:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    1932:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1933:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1934:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1935:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1936:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1937:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1938:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1939:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1940:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1941:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1942:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1943:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1944:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1945:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1946:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1947:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1948:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1949:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1950:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1951:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1952:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1953:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1954:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1955:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1956:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1957:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1958:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1959:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1960:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1961:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1962:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1963:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1964:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1965:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1966:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1967:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1968:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1969:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1970:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1971:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1972:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1973:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1974:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1975:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1976:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1977:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1978:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1979:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1980:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1981:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1982:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1983:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1984:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1985:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1986:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1987:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1988:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    1989:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1990:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1991:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1992:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    1993:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1994:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1995:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    1996:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1997:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    1998:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    1999:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2000:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2001:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2002:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2003:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2004:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2005:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2006:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2007:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2008:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2009:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2010:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2011:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2012:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2013:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2014:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2015:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2016:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2017:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2018:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2019:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2020:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2021:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2022:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2023:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2024:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2025:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2026:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2027:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2028:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2029:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2030:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2031:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2032:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2033:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2034:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2035:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2036:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2037:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2038:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2039:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2040:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2041:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2042:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2043:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2044:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2045:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2046:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2047:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2048:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2049:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2050:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2051:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2052:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 7);
    end
    2053:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2054:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2055:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2056:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2057:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2058:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2059:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2060:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2061:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2062:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2063:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2064:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2065:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2066:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2067:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2068:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2069:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2070:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2071:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2072:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2073:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2074:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2075:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2076:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2077:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2078:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2079:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2080:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2081:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2082:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2083:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2084:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2085:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2086:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2087:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2088:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2089:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2090:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2091:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2092:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2093:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2094:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2095:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2096:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2097:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2098:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2099:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2100:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2101:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2102:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2103:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2104:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2105:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2106:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2107:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2108:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2109:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2110:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2111:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2112:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2113:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2114:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2115:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2116:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2117:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2118:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2119:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2120:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2121:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2122:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2123:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2124:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2125:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2126:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2127:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2128:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2129:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2130:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2131:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2132:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2133:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2134:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2135:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2136:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2137:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2138:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2139:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2140:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2141:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2142:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2143:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2144:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2145:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2146:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2147:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2148:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2149:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2150:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2151:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2152:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2153:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2154:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2155:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2156:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2157:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2158:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2159:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2160:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2161:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2162:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2163:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2164:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2165:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2166:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2167:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2168:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2169:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2170:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2171:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2172:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2173:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2174:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2175:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2176:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2177:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2178:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2179:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2180:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2181:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2182:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2183:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2184:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2185:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2186:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2187:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2188:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2189:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2190:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2191:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2192:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2193:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2194:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2195:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2196:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2197:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2198:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2199:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2200:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2201:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2202:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2203:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2204:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2205:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2206:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2207:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2208:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2209:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2210:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2211:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2212:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2213:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2214:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2215:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2216:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2217:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2218:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2219:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2220:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2221:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2222:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2223:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2224:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2225:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2226:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2227:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2228:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2229:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2230:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2231:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2232:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2233:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2234:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2235:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2236:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2237:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2238:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2239:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2240:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2241:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2242:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2243:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2244:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2245:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2246:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2247:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2248:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2249:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2250:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2251:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2252:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2253:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2254:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2255:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2256:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2257:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2258:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2259:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2260:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2261:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2262:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2263:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2264:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2265:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2266:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2267:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2268:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2269:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2270:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2271:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2272:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2273:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2274:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2275:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2276:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2277:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2278:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2279:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2280:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2281:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2282:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2283:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2284:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2285:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2286:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2287:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2288:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2289:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2290:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2291:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2292:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2293:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2294:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2295:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2296:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2297:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2298:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2299:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2300:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2301:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2302:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2303:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2304:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2305:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2306:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2307:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2308:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2309:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2310:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2311:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2312:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2313:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2314:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2315:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2316:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2317:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2318:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2319:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2320:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2321:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2322:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2323:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2324:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2325:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2326:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2327:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2328:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2329:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2330:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2331:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2332:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2333:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2334:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2335:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2336:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2337:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2338:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2339:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2340:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2341:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2342:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2343:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2344:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2345:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2346:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2347:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2348:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2349:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2350:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2351:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2352:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2353:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2354:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2355:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2356:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2357:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2358:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2359:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2360:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2361:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2362:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2363:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2364:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2365:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2366:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2367:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2368:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2369:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2370:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2371:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2372:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2373:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2374:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2375:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2376:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2377:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2378:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2379:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2380:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2381:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2382:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2383:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2384:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2385:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2386:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2387:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2388:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2389:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2390:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2391:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2392:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2393:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2394:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2395:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2396:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2397:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2398:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2399:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2400:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2401:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2402:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2403:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2404:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2405:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2406:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2407:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2408:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2409:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2410:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2411:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2412:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2413:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2414:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2415:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2416:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2417:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2418:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2419:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2420:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2421:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2422:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2423:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2424:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2425:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2426:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2427:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2428:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2429:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2430:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2431:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2432:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2433:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2434:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2435:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2436:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2437:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2438:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2439:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2440:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2441:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2442:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2443:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2444:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2445:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2446:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2447:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2448:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2449:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2450:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2451:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2452:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2453:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2454:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2455:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2456:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2457:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2458:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2459:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2460:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2461:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2462:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2463:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2464:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2465:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2466:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2467:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2468:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2469:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2470:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2471:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2472:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2473:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2474:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2475:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2476:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2477:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2478:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2479:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2480:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2481:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2482:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2483:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2484:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2485:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2486:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2487:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2488:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2489:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2490:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2491:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2492:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2493:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2494:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2495:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2496:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2497:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2498:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2499:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2500:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2501:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2502:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2503:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2504:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2505:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2506:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2507:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2508:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2509:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2510:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2511:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2512:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2513:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2514:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2515:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2516:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2517:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2518:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2519:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2520:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2521:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2522:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2523:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2524:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2525:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2526:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2527:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2528:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2529:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2530:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2531:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2532:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2533:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2534:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2535:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2536:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2537:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2538:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2539:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2540:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2541:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2542:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2543:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2544:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2545:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2546:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2547:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2548:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2549:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2550:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2551:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2552:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2553:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2554:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2555:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2556:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2557:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2558:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2559:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2560:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2561:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2562:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2563:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2564:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2565:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2566:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2567:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2568:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2569:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2570:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2571:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2572:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2573:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2574:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2575:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2576:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2577:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2578:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2579:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2580:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2581:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2582:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2583:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2584:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2585:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2586:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2587:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2588:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2589:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2590:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2591:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2592:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2593:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2594:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2595:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2596:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2597:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2598:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2599:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2600:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2601:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2602:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2603:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2604:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2605:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2606:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2607:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2608:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2609:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 12);
    end
    2610:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2611:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2612:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2613:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2614:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2615:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2616:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2617:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2618:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2619:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2620:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2621:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2622:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2623:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2624:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2625:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2626:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2627:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2628:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2629:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2630:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2631:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2632:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2633:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2634:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2635:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2636:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2637:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2638:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2639:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2640:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2641:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2642:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2643:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2644:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2645:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2646:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2647:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2648:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2649:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2650:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2651:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2652:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2653:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2654:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2655:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2656:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2657:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2658:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2659:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2660:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2661:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2662:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2663:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2664:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2665:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2666:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2667:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2668:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2669:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2670:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2671:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2672:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 9);
    end
    2673:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2674:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2675:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 13);
    end
    2676:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2677:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2678:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2679:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2680:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2681:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2682:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2683:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2684:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2685:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2686:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2687:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2688:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2689:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2690:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2691:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2692:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2693:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2694:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2695:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2696:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2697:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2698:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2699:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2700:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2701:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2702:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2703:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2704:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2705:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2706:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2707:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 10);
    end
    2708:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2709:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2710:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2711:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2712:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2713:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2714:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2715:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2716:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2717:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2718:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2719:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2720:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2721:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2722:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2723:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2724:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2725:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2726:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2727:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2728:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2729:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2730:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2731:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2732:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2733:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2734:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2735:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2736:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2737:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2738:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2739:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2740:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2741:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2742:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2743:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2744:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2745:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2746:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2747:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2748:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2749:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2750:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2751:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2752:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2753:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2754:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2755:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2756:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2757:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2758:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2759:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2760:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2761:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2762:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2763:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2764:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2765:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2766:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2767:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2768:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2769:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2770:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2771:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2772:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2773:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2774:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2775:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2776:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2777:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2778:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2779:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2780:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2781:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2782:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2783:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2784:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2785:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2786:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2787:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2788:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2789:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2790:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2791:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2792:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2793:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2794:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2795:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2796:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2797:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2798:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2799:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2800:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2801:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2802:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2803:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2804:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2805:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2806:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2807:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2808:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2809:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2810:
    begin
        tile_x_pos = (RECT_WIDTH * 3);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2811:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2812:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2813:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2814:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2815:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2816:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2817:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2818:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2819:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2820:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2821:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2822:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2823:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2824:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2825:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2826:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2827:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2828:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2829:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2830:
    begin
        tile_x_pos = (RECT_WIDTH * 9);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2831:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2832:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2833:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2834:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2835:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2836:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2837:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2838:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2839:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2840:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2841:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2842:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2843:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2844:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2845:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2846:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2847:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2848:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2849:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2850:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2851:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2852:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2853:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2854:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2855:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2856:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2857:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2858:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2859:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2860:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2861:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2862:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2863:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2864:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2865:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2866:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2867:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2868:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2869:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2870:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2871:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2872:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2873:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2874:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2875:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2876:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2877:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2878:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2879:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2880:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2881:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2882:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2883:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2884:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2885:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2886:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2887:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2888:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2889:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2890:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2891:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2892:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2893:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2894:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2895:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2896:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 11);
    end
    2897:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2898:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2899:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2900:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2901:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2902:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2903:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2904:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2905:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2906:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2907:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2908:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2909:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2910:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2911:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2912:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2913:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2914:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2915:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2916:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2917:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2918:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2919:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2920:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2921:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2922:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2923:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2924:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2925:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2926:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2927:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2928:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2929:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2930:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2931:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2932:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2933:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2934:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2935:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 1);
    end
    2936:
    begin
        tile_x_pos = (RECT_WIDTH * 7);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2937:
    begin
        tile_x_pos = (RECT_WIDTH * 8);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2938:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2939:
    begin
        tile_x_pos = (RECT_WIDTH * 10);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2940:
    begin
        tile_x_pos = (RECT_WIDTH * 11);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2941:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2942:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 5);
    end
    2943:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2944:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2945:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2946:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2947:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2948:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2949:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2950:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2951:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2952:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2953:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2954:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2955:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2956:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    2957:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2958:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2959:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2960:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 8);
    end
    2961:
    begin
        tile_x_pos = (RECT_WIDTH * 12);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2962:
    begin
        tile_x_pos = (RECT_WIDTH * 13);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2963:
    begin
        tile_x_pos = (RECT_WIDTH * 14);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2964:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2965:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2966:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2967:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2968:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2969:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2970:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2971:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2972:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2973:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2974:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2975:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2976:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2977:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2978:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2979:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2980:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2981:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2982:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2983:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2984:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2985:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2986:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2987:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2988:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2989:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2990:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2991:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2992:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2993:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2994:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2995:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2996:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2997:
    begin
        tile_x_pos = (RECT_WIDTH * 15);
        tile_y_pos = (RECT_LENGTH * 14);
    end
    2998:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    2999:
    begin
        tile_x_pos = (RECT_WIDTH * 1);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    3000:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    3001:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3002:
    begin
        tile_x_pos = (RECT_WIDTH * 2);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3003:
    begin
        tile_x_pos = (RECT_WIDTH * 4);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    3004:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3005:
    begin
        tile_x_pos = (RECT_WIDTH * 5);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    3006:
    begin
        tile_x_pos = (RECT_WIDTH * 6);
        tile_y_pos = (RECT_LENGTH * 6);
    end
    3007:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3008:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3009:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3010:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3011:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3012:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3013:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3014:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3015:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3016:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3017:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3018:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3019:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3020:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3021:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3022:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3023:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3024:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3025:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3026:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3027:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3028:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3029:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3030:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3031:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3032:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3033:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3034:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3035:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3036:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3037:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3038:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3039:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3040:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3041:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3042:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3043:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3044:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3045:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3046:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3047:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3048:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3049:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3050:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3051:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3052:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3053:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3054:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3055:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3056:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3057:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3058:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3059:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3060:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3061:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3062:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3063:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3064:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3065:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3066:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3067:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3068:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3069:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3070:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    3071:
    begin
        tile_x_pos = (RECT_WIDTH * 0);
        tile_y_pos = (RECT_LENGTH * 0);
    end
    default:
    begin
        tile_x_pos = 0;
        tile_y_pos = 0;
    end
endcase

delay #(11, 2) hcount_delay(
 .clk(pclk),
 .rst(rst),
 .din(hcount_in),
 .dout(hcount_delayed)
);

delay #(11, 2) vcount_delay(
 .clk(pclk),
 .rst(rst),
 .din(vcount_in),
 .dout(vcount_delayed)
);

delay #(1, 2) vsync_delay(
 .clk(pclk),
 .rst(rst),
 .din(vsync_in),
 .dout(vsync_delayed)
);

delay #(1, 2) hsync_delay(
 .clk(pclk),
 .rst(rst),
 .din(hsync_in),
 .dout(hsync_delayed)
);

delay #(1, 2) vblnk_delay(
 .clk(pclk),
 .rst(rst),
 .din(vblnk_in),
 .dout(vblnk_delayed)
);

delay #(1, 2) hblnk_delay(
 .clk(pclk),
 .rst(rst),
 .din(hblnk_in),
 .dout(hblnk_delayed)
);

endmodule
